`define DATA_ADDR_BUS 31:0
`define DATA_BUS 31:0
`define DATA_MEM_NUM 131071
`define DATA_ADDR_BUS_WIDTH 17
`define BYTE_WIDTH 7:0