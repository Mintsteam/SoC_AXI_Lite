//CP0�Ĵ�����ַ
`define CP0_REG_BadVAddr    5'b01000        //ֻ��
`define CP0_REG_COUNT    5'b01001        //�ɶ�д
`define CP0_REG_COMPARE    5'b01011      //�ɶ�д
`define CP0_REG_STATUS    5'b01100       //�ɶ�д
`define CP0_REG_CAUSE    5'b01101        //ֻ��
`define CP0_REG_EPC    5'b01110          //�ɶ�д
`define CP0_REG_PRId    5'b01111         //ֻ��
`define CP0_REG_CONFIG    5'b10000       //ֻ��